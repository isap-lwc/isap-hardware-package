../../../LWC_rtl/LWC_2pass.vhd
../../LWC_tb/LWC_TB_2pass_uut.vhd